module S_counter(clk,S_in,Mov_s,valid_s);

input       S_in;
output      valid_s
output      Mov_s;
always@(*)begin
  
end

always@(posedge clk)begin
  
end